`default_nettype none

module program_mem(input clk, rst, input [9:0] pc, output [31:0] instruction);
    reg [31:0] pmem [2047:0];
    initial begin 
        // fill regfile with intermed values
        pmem[1] = 32'b1000_1000_0000_0000_1100_0000_1110_0000;
        pmem[2] = 32'b1000_1000_0001_0000_1111_0000_1110_0000;
        pmem[3] = 32'b1000_1000_0010_0000_0000_0000_0000_0001;
        pmem[4] = 32'b1000_1000_0011_0000_0000_0000_0000_0010;
        pmem[5] = 32'b1000_1000_0100_0000_0001_0000_0000_0000;
        pmem[6] = 32'b1000_1000_0101_0000_0000_0000_0000_0100;
        pmem[7] = 32'b1000_1000_0110_0000_0000_0000_0000_0000;
        pmem[8] = 32'b1000_1000_0111_0000_1111_0010_0010_0000;
        pmem[9] = 32'b1000_1000_1000_0000_0000_0000_0010_0000;
        pmem[10] = 32'b1000_1000_1001_0000_1000_0000_0010_0001;
        pmem[11] = 32'b1000_1000_1010_0000_0000_0000_0000_0111;
        pmem[12] = 32'b1000_1000_1011_0000_0000_1000_1110_0001;
        pmem[13] = 32'b1000_1000_1100_0000_1100_0000_1111_1111;
        pmem[14] = 32'b1000_1000_1101_0000_1100_0000_1000_1000;
        pmem[15] = 32'b1000_1000_1110_0000_1100_0001_1000_1110;
        pmem[16] = 32'b1000_1000_1111_0000_1100_0011_1110_0000;

        // instr     op  alu_op i operA   operB
        pmem[17] = 32'b0001_0001_0000_1000_0001_0000_0000_0000;
        // instr     op  alu_op i operA   intermed
        pmem[18] = 32'b0001_0001_1000_1000_0001_0000_0000_1000;
        // instr     op  mem_we w_addr    data_in
        pmem[19] = 32'b0010_1000_1000_1000_0000_1111_0000_1000;
        // instr     op  mem_we r_addr    
        pmem[20] = 32'b0010_0001_1000_1000_1100_0000_0000_0000;
        // instr      op  alu_op i operA   intermed 
        pmem[21] = 32'b0001_0110_1001_1000_1100_1110_1011_0000;

        // jump instruction
        pmem[512] = 32'b1100_0000_0000_1000_1000_0000_0000_0000;
    end
    always @(posedge clk) begin 
        if (rst) begin 
            instruction <= pmem[0];
        end
        instruction <= pmem[pc];
    end
endmodule
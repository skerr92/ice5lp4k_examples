module aes(input clk, input [15:0] data, input [15:0] cypher);

endmodule